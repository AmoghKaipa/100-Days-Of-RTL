`timescale 1ns / 1ps
// Construct the class in TB
