`timescale 1ns / 1ps




module day_17(

    );
endmodule
